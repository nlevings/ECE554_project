module controlBlock(A0,A1,LS,M,CntrlSig);
	input [4:0] A0,A1,LS,M;
	output [12:0] CntrlSig;
	
	assign CntrlSig = 13'd0;
endmodule